library verilog;
use verilog.vl_types.all;
entity dividebyFSM_vlg_vec_tst is
end dividebyFSM_vlg_vec_tst;
