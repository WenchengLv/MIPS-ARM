library verilog;
use verilog.vl_types.all;
entity priority_casez_vlg_vec_tst is
end priority_casez_vlg_vec_tst;
